package timing_parameters;

parameter BUFFER_SIZE =16;
parameter TRP = 24;
parameter TCL = 24;
parameter TRCD = 24;
parameter TCWD = 20;
parameter T_BURST = 4;
parameter BANK_GROUP_WIDTH = 2;
parameter BANK_WIDTH = 2;
parameter ROW_WIDTH = 15;

endpackage