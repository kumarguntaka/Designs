/**************************************************************************
***                                                                     *** 
***         Kumar Sai Reddy, Fall, 2023									*** 
***                                                                     *** 
*************************************************************************** 
***  Filename: design.sv    Created by Kumar Sai Reddy, 3/29/2023       ***  
***  Version                Version V0p1                                ***  
***  Status                 Tested                                      ***  
***************************************************************************/

package tw_factor_pkg;

parameter shortreal W4R[0:1]={1.00, 0.00};
parameter shortreal W4I[0:1]={0.00,-1.00};

parameter shortreal W8R[0:3]={1.00, 0.707, 0.00,-0.707};
parameter shortreal W8I[0:3]={0.00,-0.707,-1.00,-0.707};

parameter shortreal W16R[0:7]={1.0000,0.9239,0.7071,0.3827,0.0000,-0.3827,-0.7071,-0.9239};
parameter shortreal W16I[0:7]={0.0000,-0.3827,-0.7071,-0.9239,-1.0000,-0.9239,-0.7071,-0.3827};

parameter shortreal W32R[0:15]={1.0000,0.9808,0.9239,0.8315,0.7071,0.5556,0.3827,0.1951,0.0000,-0.1951,-0.3827,-0.5556,-0.7071,-0.8315,-0.9239,-0.9808};
parameter shortreal W32I[0:15]={0.0000,-0.1951,-0.3827,-0.5556,-0.7071,-0.8315,-0.9239,-0.9808,-1.0000,-0.9808,-0.9239,-0.8315,-0.7071,-0.5556,-0.3827,-0.1951};

parameter shortreal W64R[0:31]={1.0000,0.9952,0.9808,0.9569,0.9239,0.8819,0.8315,0.7730,0.7071,0.6344,0.5556,0.4714,0.3827,0.2903,0.1951,0.0980,0.0000,-0.0980,-0.1951,-0.2903,-0.3827,-0.4714,-0.5556,-0.6344,-0.7071,-0.7730,-0.8315,-0.8819,-0.9239,-0.9569,-0.9808,-0.9952};
parameter shortreal W64I[0:31]={0.0000,-0.0980,-0.1951,-0.2903,-0.3827,-0.4714,-0.5556,-0.6344,-0.7071,-0.7730,-0.8315,-0.8819,-0.9239,-0.9569,-0.9808,-0.9952,-1.0000,-0.9952,-0.9808,-0.9569,-0.9239,-0.8819,-0.8315,-0.7730,-0.7071,-0.6344,-0.5556,-0.4714,-0.3827,-0.2903,-0.1951,-0.0980};

parameter shortreal W128R[0:63]={1.0000,0.9988,0.9952,0.9892,0.9808,0.9700,0.9569,0.9415,0.9239,0.9040,0.8819,0.8577,0.8315,0.8032,0.7730,0.7410,0.7071,0.6716,0.6344,0.5957,0.5556,0.5141,0.4714,0.4276,0.3827,0.3369,0.2903,0.2430,0.1951,0.1467,0.0980,0.0491,0.0000,-0.0491,-0.0980,-0.1467,-0.1951,-0.2430,-0.2903,-0.3369,-0.3827,-0.4276,-0.4714,-0.5141,-0.5556,-0.5957,-0.6344,-0.6716,-0.7071,-0.7410,-0.7730,-0.8032,-0.8315,-0.8577,-0.8819,-0.9040,-0.9239,-0.9415,-0.9569,-0.9700,-0.9808,-0.9892,-0.9952,-0.9988};
parameter shortreal W128I[0:63]={0.0000,-0.0491,-0.0980,-0.1467,-0.1951,-0.2430,-0.2903,-0.3369,-0.3827,-0.4276,-0.4714,-0.5141,-0.5556,-0.5957,-0.6344,-0.6716,-0.7071,-0.7410,-0.7730,-0.8032,-0.8315,-0.8577,-0.8819,-0.9040,-0.9239,-0.9415,-0.9569,-0.9700,-0.9808,-0.9892,-0.9952,-0.9988,-1.0000,-0.9988,-0.9952,-0.9892,-0.9808,-0.9700,-0.9569,-0.9415,-0.9239,-0.9040,-0.8819,-0.8577,-0.8315,-0.8032,-0.7730,-0.7410,-0.7071,-0.6716,-0.6344,-0.5957,-0.5556,-0.5141,-0.4714,-0.4276,-0.3827,-0.3369,-0.2903,-0.2430,-0.1951,-0.1467,-0.0980,-0.0491};

endpackage