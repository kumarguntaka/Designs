/**************************************************************************
***                                                                     *** 
***         Kumar Sai Reddy, Spring, 2024									*** 
***                                                                     *** 
*************************************************************************** 
***  Filename: design.sv    Created by Kumar Sai Reddy,           ***  
***  Version                Version V0p1                                ***  
***  Status                 Tested                                      ***  
***************************************************************************/